module simple_systolic_array_tb();
    reg clk;
    reg rst_n;
    reg [11:0] matrix_a_in;
    reg [11:0] matrix_b_in;
    reg valid_in;
    wire [23:0] matrix_c_out;
    wire valid_out;
    simple_systolic_array dut(
        .clk(clk),
        .rst_n(rst_n),
        .matrix_a_in(matrix_a_in),
        .matrix_b_in(matrix_b_in),
        .valid_in(valid_in),
        .matrix_c_out(matrix_c_out),
        .valid_out(valid_out)
    );
    initial begin
        clk = 0;
        forever #1 clk = ~clk; 
    end
    initial begin
        rst_n = 0;
        matrix_a_in = 0;
        matrix_b_in = 0;
        valid_in = 0;
        @(negedge clk);
        rst_n = 1;
        if (matrix_c_out !== 24'b0 || valid_out !== 1'b0) begin
            $display("Test failed: Initial state not zero");
        end else begin
            $display("Initial state test passed");
        end
        valid_in = 1;
        matrix_a_in = 12'h741; 
        matrix_b_in = 12'h789;
        @(negedge clk);
        matrix_a_in = 12'h852;
        matrix_b_in = 12'h456;
        @(negedge clk);
        matrix_a_in = 12'h963;
        matrix_b_in = 12'h123;
        @(negedge clk);
        valid_in = 0;
        repeat(20) @(negedge clk);
        $stop; // Stop the simulation
    end
endmodule